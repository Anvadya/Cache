`include "MainMemory.v"

module CacheController(
    input wire [31:0] memoryAddress, // last 3 bits offset 
    input wire [7:0] writeValue,
    input wire isWrite,
    input wire clk,
    output wire [7:0] outputdata
);

integer Associativity = 2; // <-----associativity------->
integer Blocks = 32; 
integer no_of_rows; 
integer no_of_columns; 

//Variable parameters
parameter indexbit = 4; //log base 2 of rows

bool hitbit;
integer tag;
integer index;
integer offset; 
integer column;

reg [7:0] tempout;

reg [27:0] TagArray [0:7][0:3];
// reg [30-log(32/Associativity):0] TagArray [0:(32/Associativity)-1][0:Associativity-1];///////////////////////
reg [63:0] DataArray [0:7][0:3];
// reg [63:0] DataArray [0:(32/Associativity)-1][0:Associativity-1];////////////////////////////////////////////
integer frequency [0:7][0:3];
// integer frequency [0:(32/Associativity)-1][0:Associativity-1];///////////////////////////////////////////////

// Initialisation

initial begin
    no_of_rows = Blocks/Associativity;
    no_of_columns = Associativity;
    for(integer i=0;i<no_of_rows;i++) begin
        for(integer j=0;j<no_of_columns;j++) begin
            TagArray[i][j]=0;
            DataArray[i][j]=0;
            frequency[i][j]=j;
        end
    end
end

// Memory Variables

reg [31:0] Address;
reg [7:0] Data;
reg [0:0] ismemWrite;
wire [7:0] outputmem;

MainMemory m1 (.Address(Address),.Data(Data),.ismemWrite(ismemWrite),.outputmem(outputmem));

initial begin
    Address=0;
    Data=0;
    ismemWrite=0;
end

always @(posedge clk) begin
    offset = memoryAddress [2:0];
    index = memoryAddress [(indexbit+2):3];
    // index = memoryAddress [2+log(32/Associativity):3];/////////////////////////////////////////////////
    tag = memoryAddress [31:(indexbit+3)];
    // tag = memoryAddress [31:3+log(32/Associativity)];//////////////////////////////////////////////////
    hitbit = 0;
    column = 0;
    for (integer i=0;i<no_of_columns;i++) begin
        if (TagArray[index][i][(28-indexbit):0]==tag && TagArray[index][i][29-indexbit]==1) begin
            hitbit = 1;
            column = i;
        end
        // if (TagArray[index][i][28-log(32/Associativity):0]==tag && TagArray[index][i][29-log(32/Associativity)]==1) begin
        //     hitbit = 1;
        //     column = i;
        // end
    end
    if (isWrite==0 && hitbit==1) begin
        for (integer i=0;i<8;i++) begin
            tempout [i] = DataArray[index][column][8*offset+i];
        end
        for (integer i=0;i<no_of_columns;i++) begin
            if (frequency[index][i]==column) begin
                for (integer j=i;j>0;j--) frequency[index][j]=frequency[index][j-1];
                frequency[index][0]=column;
            end
        end
    end
    else if (hitbit==0) begin
        column = frequency[index][no_of_columns-1];
        if (TagArray[index][column][(30-indexbit)]) begin
            Address = memoryAddress;
            Address[31:(indexbit+3)] = TagArray[index][column][(28-indexbit):0];
            for (integer i=0;i<8;i++) begin
                for (integer j=0;j<8;j++) Data[j] = DataArray[index][column][8*i+j];
                Address[2:0]=i;
                ismemWrite=1;
                ismemWrite=0;
            end        
        end
        Address = memoryAddress;
        for (integer i=0;i<8;i++) begin
            Address[2:0]=i;
            for (integer j=0;j<8;j++) DataArray[index][column][8*i+j]=outputmem[j];
        end
        if (isWrite==0) begin
            for (integer i=0;i<8;i++) tempout[i]=DataArray[index][column][8*offset+i];
        end
        TagArray[index][column][(28-indexbit):0]=tag;
        // TagArray[index][column][28-log(32/Associativity):0]=tag;////////////////////////////////////////////////////////////
        TagArray[index][column][(29-indexbit)]=1;
        // TagArray[index][column][29-log(32/Associativity)]=1;///////////////////////////////////////////////////////////////
        for (integer j=no_of_columns-1;j>0;j--) frequency[index][j]=frequency[index][j-1];
        frequency[index][0]=column;
    end
    if (isWrite) begin
        for (integer i=0;i<8;i++) begin
            DataArray[index][column][8*offset+i] = writeValue[i];
        end 
    end 
    maintb.totalno++;
    if (hitbit) maintb.hitno++;
end

assign outputdata = tempout;

endmodule

module maintb();

    reg [31:0] memoryAddress_tb; 
    reg[7:0] writeValue_tb;
    reg isWrite_tb;
    reg clk;
    wire [7:0] outputdata_tb;
    
    integer hitno;
    integer totalno;
    
    CacheController c1 (.memoryAddress(memoryAddress_tb),.writeValue(writeValue_tb),.isWrite(isWrite_tb),.outputdata(outputdata_tb),.clk(clk));
    
    initial begin
        $dumpfile("tb.vcd");
        $dumpvars(0,maintb);
        hitno=0;
        totalno=0;
        clk=0;
        writeValue_tb=9;
        isWrite_tb=1;

            memoryAddress_tb = 32'h02001f91;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003be;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006b8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f90;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003c0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003c1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01001f9c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000005;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01001f9d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000002;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000760;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000761;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000762;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000763;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000764;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000765;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000766;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000767;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000768;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000769;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000770;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000771;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000772;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000773;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000774;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000775;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000776;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000777;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000778;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000779;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000780;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000781;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000782;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000783;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000784;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000785;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000786;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000787;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000788;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000789;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000790;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000791;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000792;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000793;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000794;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000795;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000796;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000797;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000798;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000799;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007aa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ab;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ac;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ad;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ae;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007af;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ba;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007be;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ca;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ce;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000001;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000000;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f83;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f84;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f85;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007da;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007db;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000800;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000801;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000802;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000803;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000804;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000805;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000806;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000807;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000808;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000809;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000810;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000811;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000812;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000813;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000814;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000815;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000816;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000817;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000818;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000819;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000820;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000821;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000822;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000823;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000824;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000825;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000826;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000827;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000828;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000829;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000830;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000831;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000832;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000833;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000834;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000835;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000836;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000837;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000838;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000839;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000840;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000841;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000842;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000843;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000844;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000845;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000846;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000847;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000848;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000849;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000850;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000851;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000852;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000853;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000854;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000855;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000856;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000857;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000858;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000859;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000760;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000761;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000762;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000763;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000764;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000765;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000766;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000767;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000768;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000769;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000770;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000771;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000772;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000773;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000774;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000775;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000776;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000777;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000778;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000779;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000780;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000781;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000782;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000783;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000784;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000785;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000786;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000806;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000787;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000788;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000789;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000806;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000790;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000791;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000792;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000793;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000794;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000795;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000796;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000816;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000797;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000798;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000799;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000816;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000826;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007aa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ab;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000826;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ac;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ad;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ae;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007af;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000836;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ba;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000836;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007be;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000846;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ca;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000846;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ce;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000856;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007da;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007db;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000856;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000760;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000761;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000762;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000763;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000764;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000765;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000766;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000767;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000768;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000769;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000770;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000771;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000772;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000773;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000774;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000775;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000776;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000777;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000778;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000779;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000780;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000781;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000782;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000783;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000784;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000785;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000786;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000806;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000787;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000788;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000789;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000806;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000790;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000791;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000792;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000793;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000794;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000795;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000796;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000816;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000797;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000798;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000799;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000816;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000826;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007aa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ab;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000826;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ac;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ad;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ae;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007af;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000836;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ba;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000836;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007be;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000846;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ca;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000846;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ce;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000856;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000706;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000716;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007da;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000726;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007db;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000736;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000856;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000746;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000756;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000760;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000761;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000762;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000763;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000764;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000765;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000766;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000767;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000768;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000769;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000770;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000771;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000772;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000773;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000774;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000775;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000776;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000777;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000778;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000779;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000780;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000781;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000782;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000783;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000784;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000785;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000786;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000807;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000787;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000788;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000789;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000807;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000790;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000791;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000792;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000793;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000794;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000795;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000796;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000817;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000797;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000798;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000799;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000817;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000827;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007aa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ab;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000827;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ac;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ad;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ae;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007af;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000837;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ba;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000837;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007be;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000847;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ca;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000847;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ce;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000857;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007da;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007db;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000857;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000760;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000761;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000762;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000763;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000764;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000765;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000766;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000767;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000768;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000769;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000770;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000771;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000772;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000773;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000774;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000775;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000776;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000777;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000778;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000779;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000780;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000781;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000782;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000783;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000784;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000785;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000786;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000807;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000787;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000788;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000789;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000807;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000790;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000791;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000792;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000793;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000794;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000795;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000796;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000817;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000797;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000798;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000799;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000817;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000827;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007aa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ab;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000827;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ac;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ad;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ae;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007af;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000837;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ba;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000837;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007be;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000847;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ca;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000847;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ce;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000857;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000707;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000717;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007da;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000727;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007db;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000737;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000857;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000747;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000757;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000760;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000761;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000762;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000763;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000764;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000765;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000766;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000767;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000768;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000769;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000770;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000771;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000772;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000773;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000774;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000775;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000776;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000777;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000778;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000779;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000800;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000780;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000781;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000782;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000783;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000800;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000784;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000785;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000786;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000808;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000787;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000788;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000789;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000808;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000810;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000790;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000791;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000792;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000793;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000810;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000794;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000795;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000796;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000818;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000797;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000798;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000799;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000818;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000820;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000820;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000828;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007aa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ab;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000828;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ac;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ad;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ae;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000830;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007af;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000830;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000838;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ba;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000838;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007be;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000840;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000840;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000848;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ca;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000848;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ce;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000850;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000850;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000858;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007da;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007db;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000858;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000760;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000761;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000762;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000763;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000764;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000765;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000766;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000767;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000768;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000769;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000770;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000771;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000772;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000773;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000774;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000775;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000776;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000777;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000778;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000779;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000800;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000780;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000781;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000782;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000783;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000800;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000784;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000785;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000786;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000808;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000787;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000788;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000789;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000808;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000810;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000790;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000791;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000792;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000793;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000810;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000794;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000795;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000796;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000818;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000797;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000798;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000799;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000818;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000820;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000820;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000828;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007aa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ab;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000828;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ac;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ad;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ae;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000830;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007af;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000830;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000838;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ba;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000838;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007be;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000840;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000840;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000848;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ca;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000848;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ce;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000850;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000850;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000858;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000700;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000708;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000710;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000718;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000720;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007da;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000728;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000730;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007db;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000738;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000858;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000740;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000748;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000750;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000758;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000760;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000761;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000762;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000763;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000764;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000765;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000766;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000767;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000768;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000769;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000770;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000771;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000772;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000773;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000774;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000775;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000776;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000777;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000778;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000779;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000801;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000780;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000781;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000782;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000783;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000801;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000784;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000785;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000786;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000809;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000787;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000788;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000789;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000809;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000811;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000790;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000791;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000792;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000793;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000811;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000794;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000795;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000796;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000819;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000797;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000798;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000799;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000819;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000821;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000821;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000829;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007aa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ab;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000829;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ac;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ad;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ae;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000831;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007af;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000831;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000839;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ba;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000839;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007be;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000841;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000841;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000849;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ca;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000849;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ce;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000851;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000851;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000859;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007da;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007db;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000859;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000760;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000761;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000762;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000763;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000764;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000765;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000766;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000767;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000768;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000769;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000770;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000771;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000772;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000773;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000774;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000775;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000776;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000777;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000778;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000779;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000801;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000780;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000781;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000782;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000783;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000801;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000784;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000785;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000786;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000809;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000787;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000788;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000789;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000809;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000811;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000790;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000791;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000792;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000793;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000811;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000794;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000795;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000796;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000819;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000797;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000798;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000799;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000819;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000821;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000821;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000829;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007aa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ab;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000829;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ac;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ad;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ae;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000831;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007af;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000831;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000839;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ba;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000839;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007be;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000841;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000841;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000849;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ca;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000849;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ce;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000851;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000851;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000859;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000701;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000709;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000711;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000719;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000721;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007da;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000729;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000731;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007db;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000739;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000859;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000741;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000749;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000751;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000759;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000760;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000761;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000762;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000763;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000764;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000765;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000766;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000767;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000768;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000769;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000770;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000771;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000772;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000773;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000774;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000775;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000776;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000777;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000778;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000779;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000802;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000780;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000781;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000782;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000783;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000802;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000784;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000785;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000786;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000787;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000788;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000789;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000812;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000790;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000791;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000792;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000793;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000812;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000794;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000795;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000796;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000797;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000798;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000799;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000822;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000822;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007aa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ab;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ac;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ad;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ae;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000832;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007af;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000832;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ba;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007be;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000842;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000842;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ca;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ce;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000852;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000852;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007da;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007db;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000760;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000761;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000762;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000763;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000764;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000765;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000766;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000767;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000768;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000769;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000770;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000771;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000772;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000773;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000774;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000775;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000776;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000777;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000778;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000779;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000802;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000780;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000781;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000782;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000783;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000802;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000784;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000785;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000786;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000787;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000788;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000789;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000812;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000790;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000791;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000792;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000793;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000812;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000794;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000795;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000796;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000797;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000798;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000799;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000822;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000822;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007aa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ab;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ac;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ad;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ae;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000832;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007af;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000832;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ba;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007be;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000842;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000842;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ca;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ce;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000852;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000852;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000702;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000712;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000722;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007da;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000732;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007db;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000742;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000752;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000760;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000761;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000762;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000763;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000764;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000765;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000766;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000767;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000768;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000769;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000770;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000771;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000772;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000773;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000774;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000775;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000776;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000777;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000778;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000779;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000803;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000780;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000781;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000782;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000783;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000803;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000784;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000785;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000786;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000787;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000788;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000789;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000813;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000790;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000791;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000792;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000793;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000813;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000794;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000795;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000796;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000797;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000798;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000799;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000823;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000823;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007aa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ab;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ac;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ad;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ae;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000833;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007af;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000833;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ba;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007be;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000843;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000843;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ca;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ce;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000853;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000853;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007da;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007db;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000760;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000761;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000762;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000763;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000764;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000765;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000766;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000767;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000768;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000769;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000770;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000771;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000772;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000773;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000774;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000775;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000776;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000777;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000778;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000779;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000803;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000780;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000781;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000782;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000783;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000803;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000784;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000785;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000786;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000787;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000788;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000789;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000813;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000790;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000791;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000792;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000793;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000813;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000794;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000795;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000796;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000797;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000798;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000799;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000823;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000823;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007aa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ab;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ac;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ad;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ae;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000833;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007af;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000833;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ba;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007be;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000843;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000843;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ca;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ce;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000853;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000853;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000703;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000713;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000723;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007da;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000733;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007db;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000743;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000753;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000760;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000761;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000762;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000763;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000764;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000765;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000766;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000767;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000768;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000769;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000770;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000771;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000772;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000773;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000774;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000775;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000776;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000777;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000778;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000779;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000804;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000780;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000781;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000782;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000783;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000804;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000784;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000785;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000786;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000787;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000788;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000789;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000814;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000790;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000791;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000792;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000793;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000814;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000794;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000795;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000796;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000797;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000798;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000799;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000824;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000824;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007aa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ab;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ac;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ad;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ae;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000834;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007af;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000834;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ba;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007be;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000844;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000844;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ca;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ce;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000854;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000854;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007da;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007db;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000760;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000761;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000762;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000763;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000764;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000765;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000766;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000767;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000768;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000769;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000770;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000771;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000772;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000773;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000774;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000775;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000776;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000777;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000778;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000779;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000804;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000780;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000781;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000782;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000783;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000804;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000784;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000785;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000786;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000787;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000788;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000789;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000814;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000790;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000791;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000792;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000793;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000814;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000794;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000795;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000796;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000797;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000798;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000799;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000824;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000824;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007aa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ab;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ac;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ad;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ae;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000834;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007af;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000834;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ba;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007be;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000844;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000844;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ca;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ce;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000854;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000854;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000704;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000714;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000724;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007da;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000734;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007db;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000744;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000754;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000760;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000761;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000762;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000763;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000764;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000765;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000766;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000767;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000768;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000769;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000770;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000771;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000772;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000773;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000774;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000775;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000776;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000777;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000778;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000779;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000805;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000780;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000781;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000782;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000783;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000805;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000784;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000785;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000786;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000787;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000788;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000789;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000815;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000790;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000791;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000792;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000793;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000815;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000794;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000795;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000796;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000797;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000798;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000799;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000825;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000825;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007aa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ab;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ac;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ad;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ae;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000835;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007af;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000835;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ba;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007be;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000845;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000845;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ca;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ce;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000855;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000855;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007da;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007db;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000760;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000761;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000762;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000763;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000764;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000765;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000766;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000767;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000768;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000769;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100076f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000770;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000771;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000772;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000773;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000774;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000775;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000776;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000777;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000778;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000779;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000805;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100077f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000780;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000781;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000782;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000783;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000805;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000784;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000785;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000786;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000787;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000788;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000789;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100080d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000815;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100078f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000790;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000791;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000792;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000793;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000815;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000794;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000795;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000796;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000797;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000798;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000799;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100081d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000825;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100079f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000825;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007a9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007aa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ab;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100082d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ac;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ad;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ae;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000835;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007af;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000835;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007b9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ba;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100083d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007be;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000845;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007bf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000845;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007c9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ca;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100084d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007ce;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000855;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007cf;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000855;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010006fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000705;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100070d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000715;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007d9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003bc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100071d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000725;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007da;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100072d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000735;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007db;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100073d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100085d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000745;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100074d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000755;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010007dd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100075d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000440;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000443;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000442;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100043f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000441;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003dc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003dd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f88;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f89;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f87;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003de;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003df;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003e0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003e1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003e2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003e3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003e4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003e5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003e6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003e7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003e8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003e9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003ea;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003eb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003ec;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003ed;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003ee;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003ef;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003f0;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003f1;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003f2;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003f3;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003f4;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003f5;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003f6;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003f7;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003f8;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003f9;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003fa;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003fb;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003fc;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003fd;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003fe;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h010003ff;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000400;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000401;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000402;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000403;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000404;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000405;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000406;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000407;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000408;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000409;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100040a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100040b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100040c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100040d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100040e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100040f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000410;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000411;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000412;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000413;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000414;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000415;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000416;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000417;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000418;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000419;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100041a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100041b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100041c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100041d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100041e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100041f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000420;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000421;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000422;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000423;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000424;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000425;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000426;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000427;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000428;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000429;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100042a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100042b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100042c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100042d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100042e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100042f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000430;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000431;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000432;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000433;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000434;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000435;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000436;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000437;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000438;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000439;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100043a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100043b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100043c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100043d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100043e;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h0100043f;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h01000442;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8c;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8a;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8b;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8d;
#10;
clk = ~clk;
#10;
clk = ~clk;
memoryAddress_tb = 32'h02001f8f;
        $display("Hits: %d",hitno);
        $display("Total: %d",totalno);
    end
endmodule