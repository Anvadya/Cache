`include "CacheController.v" 

module maintb();

    reg [31:0] memoryAddress_tb; 
    reg[7:0] writeValue_tb;
    reg isWrite_tb;
    reg clk;
    wire [7:0] outputdata_tb;
    
    integer hitno;
    integer totalno;
    
    CacheController c1 (.memoryAddress(memoryAddress_tb),.writeValue(writeValue_tb),.isWrite(isWrite_tb),.outputdata(outputdata_tb),.clk(clk));
    
    initial begin
        $dumpfile("tb.vcd");
        $dumpvars(0,maintb);
        hitno=0;
        totalno=0;
        clk=0;
        writeValue_tb=9;
        isWrite_tb=0;

        memoryAddress_tb = 32'h02001f86;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ad;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010006a0;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f85;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c7;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f60;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f61;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000440;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000498;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f75;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000499;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f76;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100049a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000003;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000002;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c7;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100049b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100049c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f72;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100049d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100049e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100049f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f75;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a0;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f76;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a1;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a2;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000003;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000002;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c7;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a3;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a4;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f73;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a5;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a6;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a7;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f75;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f76;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004aa;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000003;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000002;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c7;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004ac;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f69;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f68;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f67;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f66;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f73;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f72;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f65;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f63;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f62;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f61;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f64;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f1c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f27;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f1d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000599;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f72;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000599;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f72;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000599;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f72;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000599;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f72;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000599;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f73;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000599;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f73;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000599;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f73;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000599;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f73;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100059a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f3c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000070;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100006f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100006e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100059a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f84;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f82;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f80;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f81;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f7f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f7d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f7e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f7c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f7b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f7a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100043a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ca;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003cb;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003cc;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003cd;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ce;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003cf;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d0;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d1;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d2;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d3;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d4;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d5;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d6;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d7;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003da;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003db;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003dc;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003dd;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003de;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003df;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e0;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e1;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e2;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e3;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e4;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e5;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e6;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e7;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ea;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003eb;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ec;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ed;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ee;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ef;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f0;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f1;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f2;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f3;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f4;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f5;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f6;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f7;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003fa;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003fb;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003fc;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003fd;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003fe;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ff;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000400;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000401;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000402;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000403;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000404;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000405;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000406;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000407;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000408;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000409;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100040a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100040b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100040c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100040d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100040e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100040f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000410;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000411;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000412;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000413;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000414;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000415;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000416;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000417;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000418;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000419;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100041a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100041b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100041c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100041d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100041e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100041f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000420;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000421;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000422;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000423;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000424;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000425;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000426;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000427;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000428;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000429;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f81;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f7f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f80;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f82;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f84;
        $display("Hits: %d",hitno);
        $display("Total: %d",totalno);
    end
endmodule