`include "MainMemory.v"

module CacheController(
    input wire [31:0] memoryAddress, // last 3 bits offset 
    input wire [7:0] writeValue,
    input wire isWrite,
    input wire clk,
    output wire [7:0] outputdata
);

// <--------------------------------Variable Value to be changed-------------------------------------->
integer Blocks = 32; 
integer no_of_rows; 
integer no_of_columns; 

bool hitbit;
integer tag;
integer index;
integer offset; 
integer column;

reg [7:0] tempout;

reg [27:0] TagArray [0:7][0:3];
// reg [30-log(32/Associativity):0] TagArray [0:(32/Associativity)-1][0:Associativity-1];///////////////////////
reg [63:0] DataArray [0:7][0:3];
// reg [63:0] DataArray [0:(32/Associativity)-1][0:Associativity-1];////////////////////////////////////////////
integer frequency [0:7][0:3];
// integer frequency [0:(32/Associativity)-1][0:Associativity-1];///////////////////////////////////////////////


// Initialisation

initial begin
    no_of_rows = Blocks/Associativity;
    no_of_columns = Associativity;
    for(integer i=0;i<no_of_rows;i++) begin
        for(integer j=0;j<no_of_columns;j++) begin
            TagArray[i][j]=0;
            DataArray[i][j]=0;
            frequency[i][j]=j;
        end
    end
end

// Memory Variables

reg [31:0] Address;
reg [7:0] Data;
reg [0:0] ismemWrite;
wire [7:0] outputmem;

MainMemory m1 (.Address(Address),.Data(Data),.ismemWrite(ismemWrite),.outputmem(outputmem));

initial begin
    Address=0;
    Data=0;
    ismemWrite=0;
end

always @(posedge clk) begin
    offset = memoryAddress [2:0];
    index = memoryAddress [5:3];
    // index = memoryAddress [2+log(32/Associativity):3];/////////////////////////////////////////////////
    tag = memoryAddress [31:6];
    // tag = memoryAddress [31:3+log(32/Associativity)];//////////////////////////////////////////////////
    hitbit = 0;
    column = 0;
    for (integer i=0;i<no_of_columns;i++) begin
        if (TagArray[index][i][25:0]==tag && TagArray[index][i][26]==1) begin
            hitbit = 1;
            column = i;
        end
        // if (TagArray[index][i][28-log(32/Associativity):0]==tag && TagArray[index][i][29-log(32/Associativity)]==1) begin
        //     hitbit = 1;
        //     column = i;
        // end
    end
    if (isWrite==0 && hitbit==1) begin
        for (integer i=0;i<8;i++) begin
            tempout [i] = DataArray[index][column][8*offset+i];
        end
        for (integer i=0;i<no_of_columns;i++) begin
            if (frequency[index][i]==column) begin
                for (integer j=i;j>0;j--) frequency[index][j]=frequency[index][j-1];
                frequency[index][0]=column;
            end
        end
    end
    else if (hitbit==0) begin
        column = frequency[index][no_of_columns-1];
        if (TagArray[index][column][27]) begin
            Address = memoryAddress;
            Address[31:6] = TagArray[index][column][25:0];
            for (integer i=0;i<8;i++) begin
                for (integer j=0;j<8;j++) Data[j] = DataArray[index][column][8*i+j];
                Address[2:0]=i;
                ismemWrite=1;
                ismemWrite=0;
            end        
        end
        Address = memoryAddress;
        for (integer i=0;i<8;i++) begin
            Address[2:0]=i;
            for (integer j=0;j<8;j++) DataArray[index][column][8*i+j]=outputmem[j];
        end
        if (isWrite==0) begin
            for (integer i=0;i<8;i++) tempout[i]=DataArray[index][column][8*offset+i];
        end
        TagArray[index][column][25:0]=tag;
        // TagArray[index][column][28-log(32/Associativity):0]=tag;////////////////////////////////////////////////////////////
        TagArray[index][column][26]=1;
        // TagArray[index][column][29-log(32/Associativity)]=1;///////////////////////////////////////////////////////////////
        for (integer j=no_of_columns-1;j>0;j--) frequency[index][j]=frequency[index][j-1];
        frequency[index][0]=column;
    end
    if (isWrite) begin
        for (integer i=0;i<8;i++) begin
            DataArray[index][column][8*offset+i] = writeValue[i];
        end 
    end 
    maintb.totalno++;
    if (hitbit) maintb.hitno++;
end

assign outputdata = tempout;

endmodule

module maintb();

    reg [31:0] memoryAddress_tb; 
    reg[7:0] writeValue_tb;
    reg isWrite_tb;
    reg clk;
    wire [7:0] outputdata_tb;
    
    integer hitno;
    integer totalno;
    
    CacheController c1 (.memoryAddress(memoryAddress_tb),.writeValue(writeValue_tb),.isWrite(isWrite_tb),.outputdata(outputdata_tb),.clk(clk));
    
    initial begin
        $dumpfile("tb.vcd");
        $dumpvars(0,maintb);
        hitno=0;
        totalno=0;
        clk=0;
        writeValue_tb=9;
        isWrite_tb=1;
        memoryAddress_tb = 32'h02001f86;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ad;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010006a0;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f85;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c7;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f60;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f61;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000440;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000498;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f75;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000499;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f76;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100049a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000003;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000002;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c7;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100049b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100049c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f72;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100049d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100049e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100049f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f75;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a0;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f76;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a1;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a2;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000003;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000002;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c7;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a3;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a4;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f73;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a5;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a6;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a7;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f75;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f76;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004a9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004aa;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000003;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000002;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c7;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010004ac;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f69;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f68;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f67;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f66;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f73;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f72;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f65;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f63;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f62;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f61;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f64;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f1c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f27;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f1d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000599;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f72;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000599;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f72;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000599;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f72;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000599;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f72;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000599;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f73;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000599;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f73;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000599;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f73;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000599;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f73;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100059a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f43;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f30;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ab;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f51;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f50;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100008a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f70;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f4f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f3c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000070;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100006f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100006e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f53;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100059a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f29;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f2b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f6f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f74;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f71;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f84;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f82;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f80;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f81;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f7f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f7d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f7e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f7c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003c9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f7b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f7a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ae;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100043a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ca;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003cb;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003cc;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003cd;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ce;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003cf;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d0;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d1;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d2;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d3;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d4;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d5;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d6;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d7;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003d9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003da;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003db;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003dc;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003dd;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003de;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003df;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e0;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e1;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e2;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e3;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e4;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e5;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e6;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e7;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003e9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ea;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003eb;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ec;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ed;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ee;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ef;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f0;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f1;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f2;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f3;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f4;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f5;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f6;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f7;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f8;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003f9;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003fa;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003fb;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003fc;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003fd;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003fe;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h010003ff;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000400;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000401;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000402;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000403;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000404;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000405;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000406;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000407;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000408;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000409;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100040a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100040b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100040c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100040d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100040e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100040f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000410;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000411;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000412;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000413;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000414;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000415;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000416;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000417;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000418;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000419;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100041a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100041b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100041c;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100041d;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100041e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100041f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000420;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000421;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000422;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000423;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000424;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000425;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000426;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000427;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000428;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h01000429;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042a;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042b;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h0100042e;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f81;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f7f;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f80;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        memoryAddress_tb = 32'h02001f82;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        isWrite_tb=0;
        memoryAddress_tb = 32'h02001f85;
        #10;
        clk = ~clk;
        #10;
        clk = ~clk;
        $display("Hits: %d",hitno);
        $display("Total: %d",totalno);
    end
endmodule